`define BEHAVIOR
`define CYCLE 10.0
`define c2q 0.001
`timescale 1ns/1ps